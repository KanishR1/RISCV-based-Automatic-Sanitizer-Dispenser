VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper
  CLASS BLOCK ;
  FOREIGN wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 1155.025 BY 1165.745 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -11.980 -6.620 -10.380 1170.780 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.980 -6.620 1166.580 -5.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.980 1169.180 1166.580 1170.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 1164.980 -6.620 1166.580 1170.780 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.940 -13.220 32.540 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.540 -13.220 186.140 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.540 1092.480 186.140 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.140 -13.220 339.740 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.140 1093.100 339.740 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 491.740 -13.220 493.340 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 491.740 1093.100 493.340 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 645.340 -13.220 646.940 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 798.940 -13.220 800.540 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 952.540 -13.220 954.140 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1106.140 -13.220 1107.740 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 36.630 1173.180 38.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 189.810 1173.180 191.410 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 342.990 1173.180 344.590 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 496.170 1173.180 497.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 649.350 1173.180 650.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 802.530 1173.180 804.130 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 955.710 1173.180 957.310 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1108.890 1173.180 1110.490 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -18.580 -13.220 -16.980 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 -13.220 1173.180 -11.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1175.780 1173.180 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.580 -13.220 1173.180 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.540 -13.220 39.140 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.140 -13.220 192.740 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 191.140 1093.100 192.740 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.740 -13.220 346.340 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.740 1093.100 346.340 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.340 -13.220 499.940 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.340 1093.100 499.940 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 651.940 -13.220 653.540 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 805.540 -13.220 807.140 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.140 -13.220 960.740 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1112.740 -13.220 1114.340 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 43.230 1173.180 44.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 196.410 1173.180 198.010 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 349.590 1173.180 351.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 502.770 1173.180 504.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 655.950 1173.180 657.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 809.130 1173.180 810.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 962.310 1173.180 963.910 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1115.490 1173.180 1117.090 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -15.280 -9.920 -13.680 1174.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -15.280 -9.920 1169.880 -8.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -15.280 1172.480 1169.880 1174.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1168.280 -9.920 1169.880 1174.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.240 -13.220 35.840 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.840 -13.220 189.440 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.840 1093.100 189.440 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.440 -13.220 343.040 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 341.440 1092.480 343.040 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.040 -13.220 496.640 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.040 1092.480 496.640 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.640 -13.220 650.240 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 802.240 -13.220 803.840 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 955.840 -13.220 957.440 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1109.440 -13.220 1111.040 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 39.930 1173.180 41.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 193.110 1173.180 194.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 346.290 1173.180 347.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 499.470 1173.180 501.070 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 652.650 1173.180 654.250 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 805.830 1173.180 807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 959.010 1173.180 960.610 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1112.190 1173.180 1113.790 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -8.680 -3.320 -7.080 1167.480 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.680 -3.320 1163.280 -1.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -8.680 1165.880 1163.280 1167.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1161.680 -3.320 1163.280 1167.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.640 -13.220 29.240 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.240 -13.220 182.840 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 181.240 1092.480 182.840 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.840 -13.220 336.440 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.840 1093.100 336.440 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.440 -13.220 490.040 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.440 1092.480 490.040 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 642.040 -13.220 643.640 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 795.640 -13.220 797.240 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 949.240 -13.220 950.840 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1102.840 -13.220 1104.440 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 33.330 1173.180 34.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 186.510 1173.180 188.110 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 339.690 1173.180 341.290 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 492.870 1173.180 494.470 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 646.050 1173.180 647.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 799.230 1173.180 800.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 952.410 1173.180 954.010 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1105.590 1173.180 1107.190 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END clk
  PIN input_gpio_pins[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.025 387.640 1155.025 388.240 ;
    END
  END input_gpio_pins[0]
  PIN input_gpio_pins[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.025 394.440 1155.025 395.040 ;
    END
  END input_gpio_pins[1]
  PIN instructions[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END instructions[0]
  PIN instructions[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END instructions[1]
  PIN instructions[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END instructions[2]
  PIN output_gpio_pins[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.025 404.640 1155.025 405.240 ;
    END
  END output_gpio_pins[0]
  PIN output_gpio_pins[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.025 401.240 1155.025 401.840 ;
    END
  END output_gpio_pins[1]
  PIN output_gpio_pins[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1151.025 418.240 1155.025 418.840 ;
    END
  END output_gpio_pins[2]
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END resetn
  PIN uart_rx_break
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END uart_rx_break
  PIN uart_rx_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END uart_rx_data[0]
  PIN uart_rx_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END uart_rx_data[1]
  PIN uart_rx_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END uart_rx_data[2]
  PIN uart_rx_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END uart_rx_data[3]
  PIN uart_rx_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END uart_rx_data[4]
  PIN uart_rx_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END uart_rx_data[5]
  PIN uart_rx_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END uart_rx_data[6]
  PIN uart_rx_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END uart_rx_data[7]
  PIN uart_rx_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END uart_rx_en
  PIN uart_rx_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END uart_rx_valid
  PIN uart_rxd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END uart_rxd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 1160.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 1156.680 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 1159.280 1156.680 1160.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1155.080 3.280 1156.680 1160.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -13.220 22.640 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 -13.220 176.240 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 522.480 176.240 695.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 1092.480 176.240 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 -13.220 329.840 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 523.100 329.840 695.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 1093.100 329.840 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 -13.220 483.440 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 522.480 483.440 695.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 1092.480 483.440 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 -13.220 637.040 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 -13.220 790.640 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 -13.220 944.240 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 -13.220 1097.840 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 26.730 1173.180 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 179.910 1173.180 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 333.090 1173.180 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 486.270 1173.180 487.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 639.450 1173.180 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 792.630 1173.180 794.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 945.810 1173.180 947.410 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1098.990 1173.180 1100.590 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 1164.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 1159.980 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 1162.580 1159.980 1164.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.380 -0.020 1159.980 1164.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -13.220 25.940 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 -13.220 179.540 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 522.480 179.540 695.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 1092.480 179.540 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 -13.220 333.140 124.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 522.480 333.140 694.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 1093.100 333.140 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 -13.220 486.740 125.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 522.480 486.740 695.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 1093.100 486.740 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 -13.220 640.340 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 -13.220 793.940 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 -13.220 947.540 1177.380 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.540 -13.220 1101.140 1177.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 30.030 1173.180 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 183.210 1173.180 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 336.390 1173.180 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 489.570 1173.180 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 642.750 1173.180 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 795.930 1173.180 797.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 949.110 1173.180 950.710 ;
    END
    PORT
      LAYER met5 ;
        RECT -18.580 1102.290 1173.180 1103.890 ;
    END
  END vssd1
  PIN write_done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END write_done
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1149.080 1153.365 ;
      LAYER met1 ;
        RECT 0.000 0.000 1149.080 1153.520 ;
        RECT 0.000 -0.070 0.345 0.000 ;
        RECT 168.590 -0.070 168.845 0.000 ;
        RECT 179.320 -0.070 179.630 0.000 ;
        RECT 193.430 -0.070 193.675 0.000 ;
        RECT 207.335 -0.070 207.690 0.000 ;
        RECT 217.030 -0.070 217.350 0.000 ;
        RECT 223.790 -0.070 224.045 0.000 ;
        RECT 224.710 -0.070 225.065 0.000 ;
        RECT 227.470 -0.070 227.780 0.000 ;
        RECT 231.150 -0.070 231.455 0.000 ;
        RECT 232.070 -0.070 232.380 0.000 ;
        RECT 232.530 -0.070 232.990 0.000 ;
        RECT 237.590 -0.070 237.845 0.000 ;
        RECT 255.175 -0.070 255.555 0.000 ;
        RECT 267.490 -0.070 267.795 0.000 ;
        RECT 271.780 -0.070 272.090 0.000 ;
        RECT 284.970 -0.070 285.280 0.000 ;
        RECT 288.295 -0.070 288.650 0.000 ;
        RECT 290.490 -0.070 291.410 0.000 ;
        RECT 291.560 -0.070 291.870 0.000 ;
        RECT 303.935 -0.070 304.290 0.000 ;
        RECT 311.340 -0.070 311.650 0.000 ;
        RECT 312.750 -0.070 313.075 0.000 ;
        RECT 331.890 -0.070 332.245 0.000 ;
        RECT 333.730 -0.070 333.985 0.000 ;
        RECT 335.215 -0.070 335.570 0.000 ;
        RECT 336.595 -0.070 337.205 0.000 ;
        RECT 343.080 -0.070 343.390 0.000 ;
        RECT 352.695 -0.070 353.050 0.000 ;
        RECT 354.535 -0.070 354.890 0.000 ;
        RECT 363.170 -0.070 363.495 0.000 ;
        RECT 365.470 -0.070 365.930 0.000 ;
        RECT 372.370 -0.070 372.695 0.000 ;
        RECT 373.750 -0.070 374.100 0.000 ;
        RECT 381.215 -0.070 381.570 0.000 ;
        RECT 385.250 -0.070 385.565 0.000 ;
        RECT 393.175 -0.070 393.530 0.000 ;
        RECT 396.890 -0.070 397.210 0.000 ;
        RECT 405.595 -0.070 406.205 0.000 ;
        RECT 406.410 -0.070 406.735 0.000 ;
        RECT 411.470 -0.070 411.825 0.000 ;
        RECT 416.175 -0.070 416.530 0.000 ;
        RECT 418.370 -0.070 418.690 0.000 ;
        RECT 419.290 -0.070 419.630 0.000 ;
        RECT 428.490 -0.070 428.845 0.000 ;
        RECT 429.410 -0.070 429.665 0.000 ;
        RECT 429.870 -0.070 430.195 0.000 ;
        RECT 434.930 -0.070 435.185 0.000 ;
        RECT 439.655 -0.070 439.990 0.000 ;
        RECT 441.935 -0.070 442.750 0.000 ;
        RECT 443.670 -0.070 443.925 0.000 ;
        RECT 445.660 -0.070 445.970 0.000 ;
        RECT 448.730 -0.070 449.085 0.000 ;
        RECT 449.650 -0.070 450.110 0.000 ;
        RECT 451.030 -0.070 451.355 0.000 ;
        RECT 455.780 -0.070 456.090 0.000 ;
        RECT 457.575 -0.070 457.930 0.000 ;
        RECT 458.390 -0.070 458.735 0.000 ;
        RECT 464.370 -0.070 464.625 0.000 ;
        RECT 470.915 -0.070 471.270 0.000 ;
        RECT 483.230 -0.070 483.550 0.000 ;
        RECT 485.070 -0.070 485.530 0.000 ;
        RECT 489.210 -0.070 489.670 0.000 ;
        RECT 501.170 -0.070 501.425 0.000 ;
        RECT 504.035 -0.070 504.850 0.000 ;
        RECT 507.610 -0.070 507.955 0.000 ;
        RECT 512.820 -0.070 513.130 0.000 ;
        RECT 526.470 -0.070 526.820 0.000 ;
        RECT 528.875 -0.070 529.230 0.000 ;
        RECT 531.530 -0.070 531.990 0.000 ;
        RECT 533.830 -0.070 534.145 0.000 ;
        RECT 534.750 -0.070 535.065 0.000 ;
        RECT 535.670 -0.070 535.985 0.000 ;
        RECT 538.430 -0.070 538.685 0.000 ;
        RECT 538.995 -0.070 539.605 0.000 ;
        RECT 543.030 -0.070 543.385 0.000 ;
        RECT 545.100 -0.070 545.355 0.000 ;
        RECT 545.435 -0.070 546.045 0.000 ;
        RECT 546.250 -0.070 546.605 0.000 ;
        RECT 547.630 -0.070 547.885 0.000 ;
        RECT 548.240 -0.070 548.550 0.000 ;
        RECT 556.520 -0.070 556.830 0.000 ;
        RECT 558.210 -0.070 558.465 0.000 ;
        RECT 568.440 -0.070 568.790 0.000 ;
        RECT 571.090 -0.070 571.445 0.000 ;
        RECT 572.575 -0.070 572.930 0.000 ;
        RECT 580.855 -0.070 581.465 0.000 ;
        RECT 583.050 -0.070 583.395 0.000 ;
        RECT 585.810 -0.070 586.065 0.000 ;
        RECT 586.865 -0.070 587.190 0.000 ;
        RECT 600.070 -0.070 600.420 0.000 ;
        RECT 610.650 -0.070 611.000 0.000 ;
        RECT 615.250 -0.070 615.505 0.000 ;
        RECT 617.550 -0.070 617.805 0.000 ;
        RECT 618.160 -0.070 618.470 0.000 ;
        RECT 620.000 -0.070 620.565 0.000 ;
        RECT 620.920 -0.070 621.230 0.000 ;
        RECT 629.510 -0.070 629.855 0.000 ;
        RECT 631.455 -0.070 631.810 0.000 ;
        RECT 635.135 -0.070 635.745 0.000 ;
        RECT 637.790 -0.070 638.045 0.000 ;
        RECT 641.010 -0.070 641.265 0.000 ;
        RECT 641.575 -0.070 641.955 0.000 ;
        RECT 645.715 -0.070 646.070 0.000 ;
        RECT 646.990 -0.070 647.245 0.000 ;
        RECT 651.245 -0.070 651.590 0.000 ;
        RECT 660.940 -0.070 661.250 0.000 ;
        RECT 664.050 -0.070 664.365 0.000 ;
        RECT 668.610 -0.070 668.925 0.000 ;
        RECT 676.295 -0.070 676.430 0.000 ;
        RECT 676.570 -0.070 676.890 0.000 ;
        RECT 677.350 -0.070 677.605 0.000 ;
        RECT 680.110 -0.070 680.430 0.000 ;
        RECT 681.030 -0.070 681.285 0.000 ;
        RECT 686.550 -0.070 686.865 0.000 ;
        RECT 687.010 -0.070 687.335 0.000 ;
        RECT 689.875 -0.070 690.255 0.000 ;
        RECT 690.335 -0.070 690.690 0.000 ;
        RECT 692.530 -0.070 692.785 0.000 ;
        RECT 693.555 -0.070 694.235 0.000 ;
        RECT 694.370 -0.070 694.680 0.000 ;
        RECT 695.440 -0.070 695.750 0.000 ;
        RECT 695.900 -0.070 696.210 0.000 ;
        RECT 697.280 -0.070 697.590 0.000 ;
        RECT 697.740 -0.070 698.050 0.000 ;
        RECT 699.890 -0.070 700.145 0.000 ;
        RECT 701.270 -0.070 701.525 0.000 ;
        RECT 701.880 -0.070 702.190 0.000 ;
        RECT 705.560 -0.070 705.870 0.000 ;
        RECT 707.860 -0.070 708.170 0.000 ;
        RECT 709.550 -0.070 709.860 0.000 ;
        RECT 711.035 -0.070 711.390 0.000 ;
        RECT 711.850 -0.070 712.160 0.000 ;
        RECT 714.150 -0.070 714.405 0.000 ;
        RECT 714.760 -0.070 715.070 0.000 ;
        RECT 716.140 -0.070 716.450 0.000 ;
        RECT 716.600 -0.070 716.910 0.000 ;
        RECT 717.980 -0.070 718.290 0.000 ;
        RECT 721.650 -0.070 722.225 0.000 ;
        RECT 723.810 -0.070 724.270 0.000 ;
        RECT 724.835 -0.070 725.445 0.000 ;
        RECT 726.570 -0.070 726.825 0.000 ;
        RECT 727.950 -0.070 728.260 0.000 ;
        RECT 728.975 -0.070 729.330 0.000 ;
        RECT 729.435 -0.070 729.790 0.000 ;
        RECT 732.090 -0.070 732.445 0.000 ;
        RECT 733.010 -0.070 733.265 0.000 ;
        RECT 735.770 -0.070 736.095 0.000 ;
        RECT 736.885 -0.070 737.195 0.000 ;
        RECT 738.530 -0.070 738.785 0.000 ;
        RECT 739.450 -0.070 739.705 0.000 ;
        RECT 741.395 -0.070 741.750 0.000 ;
        RECT 742.315 -0.070 742.670 0.000 ;
        RECT 742.775 -0.070 743.130 0.000 ;
        RECT 743.725 -0.070 744.050 0.000 ;
        RECT 746.350 -0.070 746.605 0.000 ;
        RECT 746.810 -0.070 747.120 0.000 ;
        RECT 749.110 -0.070 749.420 0.000 ;
        RECT 750.640 -0.070 750.950 0.000 ;
        RECT 755.550 -0.070 756.010 0.000 ;
        RECT 757.850 -0.070 758.105 0.000 ;
        RECT 758.310 -0.070 758.635 0.000 ;
        RECT 758.875 -0.070 759.230 0.000 ;
        RECT 759.690 -0.070 760.150 0.000 ;
        RECT 766.235 -0.070 766.590 0.000 ;
        RECT 767.155 -0.070 767.510 0.000 ;
        RECT 768.120 -0.070 768.430 0.000 ;
        RECT 768.580 -0.070 768.890 0.000 ;
        RECT 770.420 -0.070 770.730 0.000 ;
        RECT 773.180 -0.070 773.490 0.000 ;
        RECT 773.595 -0.070 774.410 0.000 ;
        RECT 774.515 -0.070 775.225 0.000 ;
        RECT 776.815 -0.070 777.170 0.000 ;
        RECT 779.930 -0.070 780.185 0.000 ;
        RECT 781.415 -0.070 782.025 0.000 ;
        RECT 782.230 -0.070 782.545 0.000 ;
        RECT 787.290 -0.070 787.545 0.000 ;
        RECT 788.315 -0.070 788.670 0.000 ;
        RECT 789.590 -0.070 789.900 0.000 ;
        RECT 790.970 -0.070 791.225 0.000 ;
        RECT 791.995 -0.070 792.350 0.000 ;
        RECT 792.915 -0.070 793.270 0.000 ;
        RECT 794.650 -0.070 794.905 0.000 ;
        RECT 796.640 -0.070 796.950 0.000 ;
        RECT 797.100 -0.070 797.440 0.000 ;
        RECT 801.550 -0.070 801.860 0.000 ;
        RECT 802.165 -0.070 802.470 0.000 ;
        RECT 804.415 -0.070 804.770 0.000 ;
        RECT 805.335 -0.070 805.690 0.000 ;
        RECT 805.840 -0.070 806.150 0.000 ;
        RECT 810.855 -0.070 811.530 0.000 ;
        RECT 815.350 -0.070 815.675 0.000 ;
        RECT 817.755 -0.070 818.110 0.000 ;
        RECT 819.210 -0.070 819.535 0.000 ;
        RECT 820.975 -0.070 821.585 0.000 ;
        RECT 822.710 -0.070 823.170 0.000 ;
        RECT 823.295 -0.070 823.630 0.000 ;
        RECT 824.240 -0.070 824.775 0.000 ;
        RECT 824.780 -0.070 825.035 0.000 ;
        RECT 828.690 -0.070 829.000 0.000 ;
        RECT 831.095 -0.070 831.450 0.000 ;
        RECT 832.370 -0.070 832.625 0.000 ;
        RECT 832.980 -0.070 833.290 0.000 ;
        RECT 833.750 -0.070 834.210 0.000 ;
        RECT 834.565 -0.070 835.130 0.000 ;
        RECT 835.590 -0.070 835.945 0.000 ;
        RECT 836.650 -0.070 836.970 0.000 ;
        RECT 837.110 -0.070 837.890 0.000 ;
        RECT 838.350 -0.070 838.605 0.000 ;
        RECT 843.055 -0.070 843.410 0.000 ;
        RECT 843.975 -0.070 844.330 0.000 ;
        RECT 846.320 -0.070 846.630 0.000 ;
        RECT 852.610 -0.070 852.930 0.000 ;
        RECT 855.985 -0.070 856.600 0.000 ;
        RECT 857.210 -0.070 857.520 0.000 ;
        RECT 859.050 -0.070 859.360 0.000 ;
        RECT 861.500 -0.070 862.730 0.000 ;
        RECT 864.570 -0.070 864.925 0.000 ;
        RECT 865.640 -0.070 866.260 0.000 ;
        RECT 867.790 -0.070 868.045 0.000 ;
        RECT 869.630 -0.070 870.090 0.000 ;
        RECT 870.195 -0.070 870.550 0.000 ;
        RECT 871.115 -0.070 871.470 0.000 ;
        RECT 872.035 -0.070 872.715 0.000 ;
        RECT 875.150 -0.070 875.465 0.000 ;
        RECT 876.220 -0.070 877.345 0.000 ;
        RECT 877.450 -0.070 877.705 0.000 ;
        RECT 878.370 -0.070 878.625 0.000 ;
        RECT 879.750 -0.070 880.465 0.000 ;
        RECT 881.130 -0.070 881.440 0.000 ;
        RECT 882.970 -0.070 883.325 0.000 ;
        RECT 883.430 -0.070 883.730 0.000 ;
        RECT 884.350 -0.070 884.705 0.000 ;
        RECT 884.810 -0.070 885.270 0.000 ;
        RECT 885.730 -0.070 885.985 0.000 ;
        RECT 886.650 -0.070 887.005 0.000 ;
        RECT 887.570 -0.070 887.825 0.000 ;
        RECT 888.640 -0.070 888.950 0.000 ;
        RECT 890.330 -0.070 890.585 0.000 ;
        RECT 891.250 -0.070 891.815 0.000 ;
        RECT 895.265 -0.070 895.620 0.000 ;
        RECT 895.880 -0.070 896.205 0.000 ;
        RECT 901.475 -0.070 901.830 0.000 ;
        RECT 902.290 -0.070 902.615 0.000 ;
        RECT 902.855 -0.070 903.465 0.000 ;
        RECT 903.775 -0.070 904.130 0.000 ;
        RECT 908.420 -0.070 909.040 0.000 ;
        RECT 911.135 -0.070 911.490 0.000 ;
        RECT 911.950 -0.070 912.205 0.000 ;
        RECT 915.275 -0.070 915.630 0.000 ;
        RECT 916.090 -0.070 916.345 0.000 ;
        RECT 916.550 -0.070 916.805 0.000 ;
        RECT 917.575 -0.070 917.930 0.000 ;
        RECT 918.530 -0.070 919.310 0.000 ;
        RECT 919.670 -0.070 920.485 0.000 ;
        RECT 921.255 -0.070 921.610 0.000 ;
        RECT 921.715 -0.070 922.070 0.000 ;
        RECT 922.220 -0.070 922.530 0.000 ;
        RECT 922.635 -0.070 923.345 0.000 ;
        RECT 923.555 -0.070 924.165 0.000 ;
        RECT 926.315 -0.070 926.670 0.000 ;
        RECT 928.510 -0.070 928.765 0.000 ;
        RECT 929.430 -0.070 929.745 0.000 ;
        RECT 930.500 -0.070 930.810 0.000 ;
        RECT 931.375 -0.070 931.755 0.000 ;
        RECT 931.835 -0.070 932.545 0.000 ;
        RECT 933.570 -0.070 933.925 0.000 ;
        RECT 934.030 -0.070 934.355 0.000 ;
        RECT 934.950 -0.070 935.205 0.000 ;
        RECT 935.515 -0.070 935.870 0.000 ;
        RECT 936.330 -0.070 936.645 0.000 ;
        RECT 937.250 -0.070 937.505 0.000 ;
        RECT 937.815 -0.070 938.170 0.000 ;
        RECT 939.090 -0.070 939.400 0.000 ;
        RECT 939.550 -0.070 939.895 0.000 ;
        RECT 940.010 -0.070 940.265 0.000 ;
        RECT 940.930 -0.070 941.245 0.000 ;
        RECT 943.690 -0.070 944.000 0.000 ;
        RECT 945.530 -0.070 945.990 0.000 ;
        RECT 946.450 -0.070 946.765 0.000 ;
        RECT 947.830 -0.070 948.085 0.000 ;
        RECT 951.970 -0.070 952.280 0.000 ;
        RECT 953.350 -0.070 953.660 0.000 ;
        RECT 954.270 -0.070 954.580 0.000 ;
        RECT 956.110 -0.070 956.420 0.000 ;
        RECT 956.720 -0.070 957.030 0.000 ;
        RECT 960.250 -0.070 960.575 0.000 ;
        RECT 964.850 -0.070 965.160 0.000 ;
        RECT 965.310 -0.070 965.565 0.000 ;
        RECT 966.840 -0.070 967.405 0.000 ;
        RECT 968.070 -0.070 968.990 0.000 ;
        RECT 969.140 -0.070 969.450 0.000 ;
        RECT 970.015 -0.070 970.725 0.000 ;
        RECT 972.775 -0.070 973.130 0.000 ;
        RECT 973.280 -0.070 973.845 0.000 ;
        RECT 974.155 -0.070 974.510 0.000 ;
        RECT 975.075 -0.070 975.430 0.000 ;
        RECT 975.995 -0.070 976.350 0.000 ;
        RECT 977.730 -0.070 978.535 0.000 ;
        RECT 980.135 -0.070 980.950 0.000 ;
        RECT 981.055 -0.070 981.410 0.000 ;
        RECT 983.285 -0.070 983.610 0.000 ;
        RECT 984.170 -0.070 985.090 0.000 ;
        RECT 985.240 -0.070 985.860 0.000 ;
        RECT 986.620 -0.070 986.930 0.000 ;
        RECT 987.955 -0.070 988.890 0.000 ;
        RECT 992.910 -0.070 993.265 0.000 ;
        RECT 993.520 -0.070 993.830 0.000 ;
        RECT 993.925 -0.070 994.290 0.000 ;
        RECT 994.900 -0.070 995.210 0.000 ;
        RECT 996.695 -0.070 997.050 0.000 ;
        RECT 998.535 -0.070 998.890 0.000 ;
        RECT 1001.170 -0.070 1001.495 0.000 ;
        RECT 1002.215 -0.070 1002.570 0.000 ;
        RECT 1005.195 -0.070 1005.560 0.000 ;
        RECT 1006.815 -0.070 1007.170 0.000 ;
        RECT 1008.090 -0.070 1008.400 0.000 ;
        RECT 1009.610 -0.070 1010.185 0.000 ;
        RECT 1011.310 -0.070 1011.620 0.000 ;
        RECT 1012.335 -0.070 1012.690 0.000 ;
        RECT 1012.795 -0.070 1013.150 0.000 ;
        RECT 1013.715 -0.070 1014.070 0.000 ;
        RECT 1014.175 -0.070 1014.990 0.000 ;
        RECT 1015.095 -0.070 1015.450 0.000 ;
        RECT 1015.455 -0.070 1016.220 0.000 ;
        RECT 1016.935 -0.070 1017.290 0.000 ;
        RECT 1018.350 -0.070 1019.025 0.000 ;
        RECT 1019.280 -0.070 1019.845 0.000 ;
        RECT 1020.970 -0.070 1021.295 0.000 ;
        RECT 1021.430 -0.070 1021.740 0.000 ;
        RECT 1022.455 -0.070 1022.810 0.000 ;
        RECT 1023.500 -0.070 1023.755 0.000 ;
        RECT 1024.190 -0.070 1024.445 0.000 ;
        RECT 1025.110 -0.070 1025.420 0.000 ;
        RECT 1026.135 -0.070 1026.695 0.000 ;
        RECT 1026.950 -0.070 1027.275 0.000 ;
        RECT 1028.330 -0.070 1028.640 0.000 ;
        RECT 1030.170 -0.070 1030.480 0.000 ;
        RECT 1032.470 -0.070 1032.780 0.000 ;
        RECT 1033.080 -0.070 1033.390 0.000 ;
        RECT 1033.850 -0.070 1034.105 0.000 ;
        RECT 1035.795 -0.070 1036.150 0.000 ;
        RECT 1037.530 -0.070 1037.840 0.000 ;
        RECT 1038.910 -0.070 1039.220 0.000 ;
        RECT 1041.820 -0.070 1042.130 0.000 ;
        RECT 1044.535 -0.070 1044.890 0.000 ;
        RECT 1045.040 -0.070 1045.350 0.000 ;
        RECT 1046.880 -0.070 1047.500 0.000 ;
        RECT 1048.110 -0.070 1048.570 0.000 ;
        RECT 1049.950 -0.070 1050.205 0.000 ;
        RECT 1053.780 -0.070 1054.395 0.000 ;
        RECT 1056.035 -0.070 1056.645 0.000 ;
        RECT 1058.335 -0.070 1058.690 0.000 ;
        RECT 1060.990 -0.070 1061.345 0.000 ;
        RECT 1061.555 -0.070 1061.910 0.000 ;
        RECT 1062.600 -0.070 1062.855 0.000 ;
        RECT 1062.985 -0.070 1063.290 0.000 ;
        RECT 1064.315 -0.070 1064.670 0.000 ;
        RECT 1064.775 -0.070 1065.130 0.000 ;
        RECT 1065.590 -0.070 1065.945 0.000 ;
        RECT 1066.050 -0.070 1066.875 0.000 ;
        RECT 1075.430 -0.070 1075.740 0.000 ;
        RECT 1075.815 -0.070 1076.170 0.000 ;
        RECT 1076.275 -0.070 1076.630 0.000 ;
        RECT 1077.090 -0.070 1077.550 0.000 ;
        RECT 1078.115 -0.070 1078.470 0.000 ;
        RECT 1079.955 -0.070 1080.310 0.000 ;
        RECT 1080.460 -0.070 1080.770 0.000 ;
        RECT 1081.840 -0.070 1082.150 0.000 ;
        RECT 1083.990 -0.070 1084.345 0.000 ;
        RECT 1084.450 -0.070 1084.775 0.000 ;
        RECT 1085.830 -0.070 1086.545 0.000 ;
        RECT 1088.235 -0.070 1088.900 0.000 ;
        RECT 1089.195 -0.070 1089.970 0.000 ;
        RECT 1092.420 -0.070 1092.730 0.000 ;
        RECT 1093.755 -0.070 1094.110 0.000 ;
        RECT 1100.090 -0.070 1100.400 0.000 ;
        RECT 1102.080 -0.070 1102.390 0.000 ;
        RECT 1102.540 -0.070 1102.850 0.000 ;
        RECT 1103.460 -0.070 1103.770 0.000 ;
        RECT 1104.230 -0.070 1104.585 0.000 ;
        RECT 1104.795 -0.070 1105.150 0.000 ;
        RECT 1106.175 -0.070 1106.840 0.000 ;
        RECT 1108.475 -0.070 1109.085 0.000 ;
        RECT 1111.950 -0.070 1112.275 0.000 ;
        RECT 1112.615 -0.070 1113.430 0.000 ;
        RECT 1113.890 -0.070 1115.270 0.000 ;
        RECT 1123.550 -0.070 1123.875 0.000 ;
        RECT 1124.470 -0.070 1125.285 0.000 ;
        RECT 1127.230 -0.070 1127.585 0.000 ;
        RECT 1130.095 -0.070 1130.705 0.000 ;
        RECT 1131.015 -0.070 1131.370 0.000 ;
        RECT 1134.130 -0.070 1134.475 0.000 ;
        RECT 1136.075 -0.070 1136.685 0.000 ;
        RECT 1136.890 -0.070 1137.200 0.000 ;
        RECT 1141.490 -0.070 1141.800 0.000 ;
        RECT 1141.950 -0.070 1142.260 0.000 ;
      LAYER met2 ;
        RECT 125.620 125.620 604.160 1091.880 ;
      LAYER met3 ;
        RECT 125.000 0.000 1130.840 1091.880 ;
        RECT 153.910 -0.150 154.430 0.000 ;
        RECT 192.830 -0.150 193.430 0.000 ;
        RECT 207.350 -0.150 207.690 0.000 ;
        RECT 208.150 -0.150 208.540 0.000 ;
        RECT 209.070 -0.150 209.450 0.000 ;
        RECT 213.790 -0.150 214.270 0.000 ;
        RECT 220.490 -0.150 221.070 0.000 ;
        RECT 226.090 -0.150 226.450 0.000 ;
        RECT 234.830 -0.150 235.230 0.000 ;
        RECT 244.790 -0.150 245.410 0.000 ;
        RECT 250.700 -0.150 251.090 0.000 ;
        RECT 266.410 -0.150 267.030 0.000 ;
        RECT 267.865 -0.150 268.255 0.000 ;
        RECT 271.700 -0.150 272.090 0.000 ;
        RECT 297.920 -0.150 298.310 0.000 ;
        RECT 300.065 -0.150 300.455 0.000 ;
        RECT 302.050 -0.150 302.670 0.000 ;
        RECT 307.510 -0.150 307.900 0.000 ;
        RECT 308.890 -0.150 309.280 0.000 ;
        RECT 329.590 -0.150 329.980 0.000 ;
        RECT 331.520 -0.150 331.910 0.000 ;
        RECT 336.330 -0.150 336.950 0.000 ;
        RECT 337.410 -0.150 337.970 0.000 ;
        RECT 352.430 -0.150 353.050 0.000 ;
        RECT 361.400 -0.150 361.790 0.000 ;
        RECT 364.150 -0.150 364.550 0.000 ;
        RECT 369.150 -0.150 369.540 0.000 ;
        RECT 371.350 -0.150 371.910 0.000 ;
        RECT 376.120 -0.150 376.900 0.000 ;
        RECT 378.880 -0.150 379.270 0.000 ;
        RECT 379.500 -0.150 380.020 0.000 ;
        RECT 386.010 -0.150 386.630 0.000 ;
        RECT 386.700 -0.150 387.090 0.000 ;
        RECT 387.390 -0.150 388.010 0.000 ;
        RECT 407.790 -0.150 408.180 0.000 ;
        RECT 410.465 -0.150 410.855 0.000 ;
        RECT 428.790 -0.150 429.410 0.000 ;
        RECT 433.520 -0.150 433.910 0.000 ;
        RECT 436.225 -0.150 436.615 0.000 ;
        RECT 442.130 -0.150 442.750 0.000 ;
        RECT 452.940 -0.150 453.330 0.000 ;
        RECT 455.700 -0.150 456.090 0.000 ;
        RECT 457.310 -0.150 457.930 0.000 ;
        RECT 460.990 -0.150 462.070 0.000 ;
        RECT 470.350 -0.150 470.740 0.000 ;
        RECT 484.150 -0.150 484.540 0.000 ;
        RECT 487.440 -0.150 488.220 0.000 ;
        RECT 492.040 -0.150 492.660 0.000 ;
        RECT 502.390 -0.150 503.010 0.000 ;
        RECT 504.390 -0.150 504.990 0.000 ;
        RECT 508.650 -0.150 509.840 0.000 ;
        RECT 516.880 -0.150 517.500 0.000 ;
        RECT 522.790 -0.150 523.390 0.000 ;
        RECT 524.930 -0.150 525.550 0.000 ;
        RECT 534.690 -0.150 535.210 0.000 ;
        RECT 538.430 -0.150 539.350 0.000 ;
        RECT 540.570 -0.150 541.580 0.000 ;
        RECT 545.100 -0.150 545.490 0.000 ;
        RECT 550.690 -0.150 551.310 0.000 ;
        RECT 575.070 -0.150 575.690 0.000 ;
        RECT 578.450 -0.150 578.840 0.000 ;
        RECT 610.650 -0.150 611.040 0.000 ;
        RECT 611.640 -0.150 612.260 0.000 ;
        RECT 617.780 -0.150 618.170 0.000 ;
        RECT 618.700 -0.150 619.090 0.000 ;
        RECT 620.310 -0.150 620.700 0.000 ;
        RECT 621.300 -0.150 621.690 0.000 ;
        RECT 621.760 -0.150 622.150 0.000 ;
        RECT 622.910 -0.150 623.530 0.000 ;
        RECT 624.060 -0.150 624.450 0.000 ;
        RECT 628.590 -0.150 629.110 0.000 ;
        RECT 629.350 -0.150 629.740 0.000 ;
        RECT 630.270 -0.150 630.660 0.000 ;
        RECT 630.960 -0.150 631.740 0.000 ;
        RECT 632.270 -0.150 632.660 0.000 ;
        RECT 633.260 -0.150 633.650 0.000 ;
        RECT 638.850 -0.150 639.170 0.000 ;
        RECT 639.930 -0.150 640.550 0.000 ;
        RECT 642.920 -0.150 643.310 0.000 ;
        RECT 645.610 -0.150 646.530 0.000 ;
        RECT 654.140 -0.150 654.580 0.000 ;
        RECT 656.260 -0.150 656.650 0.000 ;
        RECT 657.870 -0.150 658.490 0.000 ;
        RECT 660.400 -0.150 660.790 0.000 ;
        RECT 664.470 -0.150 665.010 0.000 ;
        RECT 665.460 -0.150 666.310 0.000 ;
        RECT 669.300 -0.150 669.900 0.000 ;
        RECT 669.990 -0.150 670.910 0.000 ;
        RECT 674.590 -0.150 674.980 0.000 ;
        RECT 676.270 -0.150 676.660 0.000 ;
        RECT 677.420 -0.150 677.810 0.000 ;
        RECT 677.880 -0.150 678.270 0.000 ;
        RECT 680.110 -0.150 680.500 0.000 ;
        RECT 680.640 -0.150 681.420 0.000 ;
        RECT 681.560 -0.150 682.340 0.000 ;
        RECT 682.480 -0.150 682.870 0.000 ;
        RECT 682.940 -0.150 683.720 0.000 ;
        RECT 697.890 -0.150 698.510 0.000 ;
        RECT 706.330 -0.150 706.900 0.000 ;
        RECT 709.620 -0.150 710.400 0.000 ;
        RECT 711.690 -0.150 712.310 0.000 ;
        RECT 714.680 -0.150 715.460 0.000 ;
        RECT 717.260 -0.150 717.830 0.000 ;
        RECT 718.980 -0.150 719.370 0.000 ;
        RECT 721.350 -0.150 721.970 0.000 ;
        RECT 724.800 -0.150 725.190 0.000 ;
        RECT 726.110 -0.150 726.500 0.000 ;
        RECT 727.100 -0.150 728.410 0.000 ;
        RECT 730.550 -0.150 731.170 0.000 ;
        RECT 731.700 -0.150 732.090 0.000 ;
        RECT 732.390 -0.150 733.470 0.000 ;
        RECT 734.250 -0.150 735.240 0.000 ;
        RECT 736.090 -0.150 736.690 0.000 ;
        RECT 739.290 -0.150 740.370 0.000 ;
        RECT 742.070 -0.150 742.670 0.000 ;
        RECT 743.660 -0.150 744.050 0.000 ;
        RECT 744.580 -0.150 745.430 0.000 ;
        RECT 746.350 -0.150 746.740 0.000 ;
        RECT 747.130 -0.150 747.730 0.000 ;
        RECT 750.100 -0.150 750.490 0.000 ;
        RECT 751.480 -0.150 751.870 0.000 ;
        RECT 753.020 -0.150 753.410 0.000 ;
        RECT 761.070 -0.150 761.460 0.000 ;
        RECT 770.800 -0.150 771.190 0.000 ;
        RECT 772.800 -0.150 773.490 0.000 ;
        RECT 774.020 -0.150 774.800 0.000 ;
        RECT 775.860 -0.150 776.250 0.000 ;
        RECT 779.770 -0.150 780.390 0.000 ;
        RECT 782.460 -0.150 783.150 0.000 ;
        RECT 783.450 -0.150 784.530 0.000 ;
        RECT 784.600 -0.150 785.450 0.000 ;
        RECT 788.740 -0.150 789.520 0.000 ;
        RECT 791.890 -0.150 792.280 0.000 ;
        RECT 798.330 -0.150 798.720 0.000 ;
        RECT 813.970 -0.150 814.360 0.000 ;
        RECT 815.880 -0.150 816.270 0.000 ;
        RECT 818.460 -0.150 819.030 0.000 ;
        RECT 819.100 -0.150 819.490 0.000 ;
        RECT 820.250 -0.150 821.330 0.000 ;
        RECT 821.650 -0.150 822.250 0.000 ;
        RECT 824.160 -0.150 825.170 0.000 ;
        RECT 827.310 -0.150 827.700 0.000 ;
        RECT 831.060 -0.150 831.450 0.000 ;
        RECT 834.530 -0.150 835.130 0.000 ;
        RECT 839.730 -0.150 840.120 0.000 ;
        RECT 845.940 -0.150 846.330 0.000 ;
        RECT 847.090 -0.150 848.010 0.000 ;
        RECT 851.760 -0.150 852.540 0.000 ;
        RECT 856.820 -0.150 857.210 0.000 ;
        RECT 857.280 -0.150 858.060 0.000 ;
        RECT 858.660 -0.150 859.050 0.000 ;
        RECT 859.580 -0.150 860.360 0.000 ;
        RECT 863.490 -0.150 864.110 0.000 ;
        RECT 868.110 -0.150 869.630 0.000 ;
        RECT 869.700 -0.150 870.090 0.000 ;
        RECT 870.550 -0.150 871.010 0.000 ;
        RECT 871.080 -0.150 871.930 0.000 ;
        RECT 872.000 -0.150 872.850 0.000 ;
        RECT 882.580 -0.150 883.360 0.000 ;
        RECT 885.340 -0.150 886.120 0.000 ;
        RECT 886.260 -0.150 887.040 0.000 ;
        RECT 889.020 -0.150 889.410 0.000 ;
        RECT 890.100 -0.150 890.490 0.000 ;
        RECT 891.090 -0.150 891.710 0.000 ;
        RECT 891.780 -0.150 892.560 0.000 ;
        RECT 894.540 -0.150 895.320 0.000 ;
        RECT 895.620 -0.150 896.010 0.000 ;
        RECT 899.600 -0.150 899.990 0.000 ;
        RECT 900.450 -0.150 901.140 0.000 ;
        RECT 901.210 -0.150 901.830 0.000 ;
        RECT 901.900 -0.150 903.320 0.000 ;
        RECT 903.740 -0.150 904.130 0.000 ;
        RECT 911.790 -0.150 912.800 0.000 ;
        RECT 913.400 -0.150 914.180 0.000 ;
        RECT 919.170 -0.150 919.770 0.000 ;
        RECT 921.220 -0.150 921.610 0.000 ;
        RECT 922.600 -0.150 922.990 0.000 ;
        RECT 924.230 -0.150 925.450 0.000 ;
        RECT 926.510 -0.150 927.130 0.000 ;
        RECT 927.660 -0.150 928.050 0.000 ;
        RECT 928.580 -0.150 929.820 0.000 ;
        RECT 930.880 -0.150 931.890 0.000 ;
        RECT 937.570 -0.150 938.170 0.000 ;
        RECT 938.930 -0.150 940.400 0.000 ;
        RECT 959.630 -0.150 960.710 0.000 ;
        RECT 964.230 -0.150 964.850 0.000 ;
        RECT 965.610 -0.150 966.230 0.000 ;
        RECT 966.990 -0.150 968.070 0.000 ;
        RECT 968.830 -0.150 969.450 0.000 ;
        RECT 969.980 -0.150 970.760 0.000 ;
        RECT 974.120 -0.150 974.510 0.000 ;
        RECT 975.040 -0.150 976.580 0.000 ;
        RECT 977.340 -0.150 977.730 0.000 ;
        RECT 980.260 -0.150 980.650 0.000 ;
        RECT 983.020 -0.150 983.410 0.000 ;
        RECT 983.780 -0.150 984.170 0.000 ;
        RECT 985.550 -0.150 985.940 0.000 ;
        RECT 987.230 -0.150 988.540 0.000 ;
        RECT 988.610 -0.150 990.150 0.000 ;
        RECT 994.590 -0.150 995.210 0.000 ;
        RECT 1000.270 -0.150 1000.660 0.000 ;
        RECT 1000.800 -0.150 1001.190 0.000 ;
        RECT 1005.400 -0.150 1005.790 0.000 ;
        RECT 1009.540 -0.150 1010.390 0.000 ;
        RECT 1011.610 -0.150 1012.690 0.000 ;
        RECT 1012.990 -0.150 1013.610 0.000 ;
        RECT 1014.830 -0.150 1016.370 0.000 ;
        RECT 1017.150 -0.150 1018.320 0.000 ;
        RECT 1019.590 -0.150 1019.980 0.000 ;
        RECT 1021.040 -0.150 1021.430 0.000 ;
        RECT 1022.210 -0.150 1022.810 0.000 ;
        RECT 1023.500 -0.150 1024.190 0.000 ;
        RECT 1030.240 -0.150 1030.630 0.000 ;
        RECT 1033.230 -0.150 1034.240 0.000 ;
        RECT 1040.360 -0.150 1040.750 0.000 ;
        RECT 1044.270 -0.150 1044.890 0.000 ;
        RECT 1052.110 -0.150 1052.710 0.000 ;
        RECT 1056.850 -0.150 1057.240 0.000 ;
        RECT 1061.980 -0.150 1063.290 0.000 ;
        RECT 1066.050 -0.150 1066.970 0.000 ;
        RECT 1068.810 -0.150 1069.200 0.000 ;
        RECT 1069.570 -0.150 1070.190 0.000 ;
        RECT 1072.790 -0.150 1073.410 0.000 ;
        RECT 1074.400 -0.150 1075.180 0.000 ;
        RECT 1078.010 -0.150 1078.400 0.000 ;
        RECT 1085.140 -0.150 1085.530 0.000 ;
        RECT 1095.350 -0.150 1096.340 0.000 ;
        RECT 1106.370 -0.150 1106.990 0.000 ;
        RECT 1108.690 -0.150 1109.290 0.000 ;
        RECT 1113.890 -0.150 1114.810 0.000 ;
        RECT 1117.640 -0.150 1118.490 0.000 ;
        RECT 1122.470 -0.150 1123.090 0.000 ;
        RECT 1124.080 -0.150 1125.320 0.000 ;
        RECT 1126.770 -0.150 1127.160 0.000 ;
        RECT 1127.530 -0.150 1128.150 0.000 ;
        RECT 1129.830 -0.150 1130.840 0.000 ;
      LAYER met4 ;
        RECT 125.620 1092.080 174.240 1092.500 ;
        RECT 176.640 1092.080 177.540 1092.500 ;
        RECT 179.940 1092.080 180.840 1092.500 ;
        RECT 183.240 1092.080 184.140 1092.500 ;
        RECT 186.540 1092.080 341.040 1092.500 ;
        RECT 343.440 1092.080 481.440 1092.500 ;
        RECT 483.840 1092.080 488.040 1092.500 ;
        RECT 490.440 1092.080 494.640 1092.500 ;
        RECT 497.040 1092.080 635.040 1092.500 ;
        RECT 125.620 695.420 635.040 1092.080 ;
        RECT 125.620 522.080 174.240 695.420 ;
        RECT 176.640 522.080 177.540 695.420 ;
        RECT 179.940 522.700 327.840 695.420 ;
        RECT 330.240 694.800 481.440 695.420 ;
        RECT 330.240 522.700 331.140 694.800 ;
        RECT 179.940 522.080 331.140 522.700 ;
        RECT 333.540 522.080 481.440 694.800 ;
        RECT 483.840 522.080 484.740 695.420 ;
        RECT 487.140 522.080 635.040 695.420 ;
        RECT 125.620 125.420 635.040 522.080 ;
        RECT 125.620 0.000 174.240 125.420 ;
        RECT 176.640 0.000 177.540 125.420 ;
        RECT 179.940 0.000 180.840 125.420 ;
        RECT 183.240 0.000 184.140 125.420 ;
        RECT 186.540 0.000 187.440 125.420 ;
        RECT 189.840 0.000 190.740 125.420 ;
        RECT 193.140 124.800 481.440 125.420 ;
        RECT 193.140 0.000 327.840 124.800 ;
        RECT 330.240 0.000 331.140 124.800 ;
        RECT 333.540 0.000 334.440 124.800 ;
        RECT 336.840 0.000 337.740 124.800 ;
        RECT 340.140 0.000 341.040 124.800 ;
        RECT 343.440 0.000 344.340 124.800 ;
        RECT 346.740 0.000 481.440 124.800 ;
        RECT 483.840 0.000 484.740 125.420 ;
        RECT 487.140 0.000 488.040 125.420 ;
        RECT 490.440 0.000 491.340 125.420 ;
        RECT 493.740 0.000 494.640 125.420 ;
        RECT 497.040 0.000 497.940 125.420 ;
        RECT 500.340 0.000 635.040 125.420 ;
        RECT 637.440 0.000 638.340 1092.500 ;
        RECT 640.740 0.000 641.640 1092.500 ;
        RECT 644.040 0.000 644.940 1092.500 ;
        RECT 647.340 0.000 648.240 1092.500 ;
        RECT 650.640 0.000 651.540 1092.500 ;
        RECT 653.940 0.000 788.640 1092.500 ;
        RECT 791.040 0.000 791.940 1092.500 ;
        RECT 794.340 0.000 795.240 1092.500 ;
        RECT 797.640 0.000 798.540 1092.500 ;
        RECT 800.940 0.000 801.840 1092.500 ;
        RECT 804.240 0.000 805.140 1092.500 ;
        RECT 807.540 0.000 942.240 1092.500 ;
        RECT 944.640 0.000 945.540 1092.500 ;
        RECT 947.940 0.000 948.840 1092.500 ;
        RECT 951.240 0.000 952.140 1092.500 ;
        RECT 954.540 0.000 955.440 1092.500 ;
        RECT 957.840 0.000 958.740 1092.500 ;
        RECT 961.140 0.000 1095.840 1092.500 ;
        RECT 1098.240 0.000 1099.140 1092.500 ;
        RECT 1101.540 0.000 1102.440 1092.500 ;
        RECT 1104.840 0.000 1105.740 1092.500 ;
        RECT 1108.140 0.000 1109.040 1092.500 ;
        RECT 1111.440 0.000 1112.340 1092.500 ;
        RECT 1114.740 0.000 1124.620 1092.500 ;
        RECT 630.510 -0.620 630.810 0.000 ;
        RECT 633.500 -0.620 633.800 0.000 ;
        RECT 677.200 -0.620 677.500 0.000 ;
        RECT 728.260 -0.620 728.560 0.000 ;
        RECT 747.580 -0.620 747.880 0.000 ;
        RECT 771.040 -0.620 771.340 0.000 ;
        RECT 785.300 -0.620 785.600 0.000 ;
        RECT 822.100 -0.620 822.400 0.000 ;
        RECT 857.520 -0.620 857.820 0.000 ;
        RECT 859.820 -0.620 860.120 0.000 ;
        RECT 862.350 -0.620 862.650 0.000 ;
        RECT 863.960 -0.620 864.260 0.000 ;
        RECT 882.820 -0.620 883.120 0.000 ;
        RECT 889.260 -0.620 889.560 0.000 ;
        RECT 889.720 -0.620 890.020 0.000 ;
        RECT 892.020 -0.620 892.320 0.000 ;
        RECT 900.990 -0.620 901.290 0.000 ;
        RECT 901.680 -0.620 901.980 0.000 ;
        RECT 912.260 -0.620 912.560 0.000 ;
        RECT 913.640 -0.620 913.940 0.000 ;
        RECT 918.700 -0.620 919.000 0.000 ;
        RECT 1012.540 -0.620 1012.840 0.000 ;
        RECT 1015.300 -0.620 1015.600 0.000 ;
        RECT 1030.480 -0.620 1030.780 0.000 ;
        RECT 1124.320 -0.620 1124.620 0.000 ;
  END
END wrapper
END LIBRARY

