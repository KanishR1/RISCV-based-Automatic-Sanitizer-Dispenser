magic
tech sky130A
magscale 1 2
timestamp 1699989578
<< obsli1 >>
rect 1104 2159 229816 230673
<< obsm1 >>
rect 0 0 229816 230704
rect 0 -14 69 0
rect 33718 -14 33769 0
rect 35864 -14 35926 0
rect 38686 -14 38735 0
rect 41467 -14 41538 0
rect 43406 -14 43470 0
rect 44758 -14 44809 0
rect 44942 -14 45013 0
rect 45494 -14 45556 0
rect 46230 -14 46291 0
rect 46414 -14 46476 0
rect 46506 -14 46598 0
rect 47518 -14 47569 0
rect 51035 -14 51111 0
rect 53498 -14 53559 0
rect 54356 -14 54418 0
rect 56994 -14 57056 0
rect 57659 -14 57730 0
rect 58098 -14 58282 0
rect 58312 -14 58374 0
rect 60787 -14 60858 0
rect 62268 -14 62330 0
rect 62550 -14 62615 0
rect 66378 -14 66449 0
rect 66746 -14 66797 0
rect 67043 -14 67114 0
rect 67319 -14 67441 0
rect 68616 -14 68678 0
rect 70539 -14 70610 0
rect 70907 -14 70978 0
rect 72634 -14 72699 0
rect 73094 -14 73186 0
rect 74474 -14 74539 0
rect 74750 -14 74820 0
rect 76243 -14 76314 0
rect 77050 -14 77113 0
rect 78635 -14 78706 0
rect 79378 -14 79442 0
rect 81119 -14 81241 0
rect 81282 -14 81347 0
rect 82294 -14 82365 0
rect 83235 -14 83306 0
rect 83674 -14 83738 0
rect 83858 -14 83926 0
rect 85698 -14 85769 0
rect 85882 -14 85933 0
rect 85974 -14 86039 0
rect 86986 -14 87037 0
rect 87931 -14 87998 0
rect 88387 -14 88550 0
rect 88734 -14 88785 0
rect 89132 -14 89194 0
rect 89746 -14 89817 0
rect 89930 -14 90022 0
rect 90206 -14 90271 0
rect 91156 -14 91218 0
rect 91515 -14 91586 0
rect 91678 -14 91747 0
rect 92874 -14 92925 0
rect 94183 -14 94254 0
rect 96646 -14 96710 0
rect 97014 -14 97106 0
rect 97842 -14 97934 0
rect 100234 -14 100285 0
rect 100807 -14 100970 0
rect 101522 -14 101591 0
rect 102564 -14 102626 0
rect 105294 -14 105364 0
rect 105775 -14 105846 0
rect 106306 -14 106398 0
rect 106766 -14 106829 0
rect 106950 -14 107013 0
rect 107134 -14 107197 0
rect 107686 -14 107737 0
rect 107799 -14 107921 0
rect 108606 -14 108677 0
rect 109020 -14 109071 0
rect 109087 -14 109209 0
rect 109250 -14 109321 0
rect 109526 -14 109577 0
rect 109648 -14 109710 0
rect 111304 -14 111366 0
rect 111642 -14 111693 0
rect 113688 -14 113758 0
rect 114218 -14 114289 0
rect 114515 -14 114586 0
rect 116171 -14 116293 0
rect 116610 -14 116679 0
rect 117162 -14 117213 0
rect 117373 -14 117438 0
rect 120014 -14 120084 0
rect 122130 -14 122200 0
rect 123050 -14 123101 0
rect 123510 -14 123561 0
rect 123632 -14 123694 0
rect 124000 -14 124113 0
rect 124184 -14 124246 0
rect 125902 -14 125971 0
rect 126291 -14 126362 0
rect 127027 -14 127149 0
rect 127558 -14 127609 0
rect 128202 -14 128253 0
rect 128315 -14 128391 0
rect 129143 -14 129214 0
rect 129398 -14 129449 0
rect 130249 -14 130318 0
rect 132188 -14 132250 0
rect 132810 -14 132873 0
rect 133722 -14 133785 0
rect 135259 -14 135286 0
rect 135314 -14 135378 0
rect 135470 -14 135521 0
rect 136022 -14 136086 0
rect 136206 -14 136257 0
rect 137310 -14 137373 0
rect 137402 -14 137467 0
rect 137975 -14 138051 0
rect 138067 -14 138138 0
rect 138506 -14 138557 0
rect 138711 -14 138847 0
rect 138874 -14 138936 0
rect 139088 -14 139150 0
rect 139180 -14 139242 0
rect 139456 -14 139518 0
rect 139548 -14 139610 0
rect 139978 -14 140029 0
rect 140254 -14 140305 0
rect 140376 -14 140438 0
rect 141112 -14 141174 0
rect 141572 -14 141634 0
rect 141910 -14 141972 0
rect 142207 -14 142278 0
rect 142370 -14 142432 0
rect 142830 -14 142881 0
rect 142952 -14 143014 0
rect 143228 -14 143290 0
rect 143320 -14 143382 0
rect 143596 -14 143658 0
rect 144330 -14 144445 0
rect 144762 -14 144854 0
rect 144967 -14 145089 0
rect 145314 -14 145365 0
rect 145590 -14 145652 0
rect 145795 -14 145866 0
rect 145887 -14 145958 0
rect 146418 -14 146489 0
rect 146602 -14 146653 0
rect 147154 -14 147219 0
rect 147377 -14 147439 0
rect 147706 -14 147757 0
rect 147890 -14 147941 0
rect 148279 -14 148350 0
rect 148463 -14 148534 0
rect 148555 -14 148626 0
rect 148745 -14 148810 0
rect 149270 -14 149321 0
rect 149362 -14 149424 0
rect 149822 -14 149884 0
rect 150128 -14 150190 0
rect 151110 -14 151202 0
rect 151570 -14 151621 0
rect 151662 -14 151727 0
rect 151775 -14 151846 0
rect 151938 -14 152030 0
rect 153247 -14 153318 0
rect 153431 -14 153502 0
rect 153624 -14 153686 0
rect 153716 -14 153778 0
rect 154084 -14 154146 0
rect 154636 -14 154698 0
rect 154719 -14 154882 0
rect 154903 -14 155045 0
rect 155363 -14 155434 0
rect 155986 -14 156037 0
rect 156283 -14 156405 0
rect 156446 -14 156509 0
rect 157458 -14 157509 0
rect 157663 -14 157734 0
rect 157918 -14 157980 0
rect 158194 -14 158245 0
rect 158399 -14 158470 0
rect 158583 -14 158654 0
rect 158930 -14 158981 0
rect 159328 -14 159390 0
rect 159420 -14 159488 0
rect 160310 -14 160372 0
rect 160433 -14 160494 0
rect 160883 -14 160954 0
rect 161067 -14 161138 0
rect 161168 -14 161230 0
rect 162171 -14 162306 0
rect 163070 -14 163135 0
rect 163551 -14 163622 0
rect 163842 -14 163907 0
rect 164195 -14 164317 0
rect 164542 -14 164634 0
rect 164659 -14 164726 0
rect 164848 -14 164955 0
rect 164956 -14 165007 0
rect 165738 -14 165800 0
rect 166219 -14 166290 0
rect 166474 -14 166525 0
rect 166596 -14 166658 0
rect 166750 -14 166842 0
rect 166913 -14 167026 0
rect 167118 -14 167189 0
rect 167330 -14 167394 0
rect 167422 -14 167578 0
rect 167670 -14 167721 0
rect 168611 -14 168682 0
rect 168795 -14 168866 0
rect 169264 -14 169326 0
rect 170522 -14 170586 0
rect 171197 -14 171320 0
rect 171442 -14 171504 0
rect 171810 -14 171872 0
rect 172300 -14 172546 0
rect 172914 -14 172985 0
rect 173128 -14 173252 0
rect 173558 -14 173609 0
rect 173926 -14 174018 0
rect 174039 -14 174110 0
rect 174223 -14 174294 0
rect 174407 -14 174543 0
rect 175030 -14 175093 0
rect 175244 -14 175469 0
rect 175490 -14 175541 0
rect 175674 -14 175725 0
rect 175950 -14 176093 0
rect 176226 -14 176288 0
rect 176594 -14 176665 0
rect 176686 -14 176746 0
rect 176870 -14 176941 0
rect 176962 -14 177054 0
rect 177146 -14 177197 0
rect 177330 -14 177401 0
rect 177514 -14 177565 0
rect 177728 -14 177790 0
rect 178066 -14 178117 0
rect 178250 -14 178363 0
rect 179053 -14 179124 0
rect 179176 -14 179241 0
rect 180295 -14 180366 0
rect 180458 -14 180523 0
rect 180571 -14 180693 0
rect 180755 -14 180826 0
rect 181684 -14 181808 0
rect 182227 -14 182298 0
rect 182390 -14 182441 0
rect 183055 -14 183126 0
rect 183218 -14 183269 0
rect 183310 -14 183361 0
rect 183515 -14 183586 0
rect 183706 -14 183862 0
rect 183934 -14 184097 0
rect 184251 -14 184322 0
rect 184343 -14 184414 0
rect 184444 -14 184506 0
rect 184527 -14 184669 0
rect 184711 -14 184833 0
rect 185263 -14 185334 0
rect 185702 -14 185753 0
rect 185886 -14 185949 0
rect 186100 -14 186162 0
rect 186275 -14 186351 0
rect 186367 -14 186509 0
rect 186714 -14 186785 0
rect 186806 -14 186871 0
rect 186990 -14 187041 0
rect 187103 -14 187174 0
rect 187266 -14 187329 0
rect 187450 -14 187501 0
rect 187563 -14 187634 0
rect 187818 -14 187880 0
rect 187910 -14 187979 0
rect 188002 -14 188053 0
rect 188186 -14 188249 0
rect 188738 -14 188800 0
rect 189106 -14 189198 0
rect 189290 -14 189353 0
rect 189566 -14 189617 0
rect 190394 -14 190456 0
rect 190670 -14 190732 0
rect 190854 -14 190916 0
rect 191222 -14 191284 0
rect 191344 -14 191406 0
rect 192050 -14 192115 0
rect 192970 -14 193032 0
rect 193062 -14 193113 0
rect 193368 -14 193481 0
rect 193614 -14 193798 0
rect 193828 -14 193890 0
rect 194003 -14 194145 0
rect 194555 -14 194626 0
rect 194656 -14 194769 0
rect 194831 -14 194902 0
rect 195015 -14 195086 0
rect 195199 -14 195270 0
rect 195546 -14 195707 0
rect 196027 -14 196190 0
rect 196211 -14 196282 0
rect 196657 -14 196722 0
rect 196834 -14 197018 0
rect 197048 -14 197172 0
rect 197324 -14 197386 0
rect 197591 -14 197778 0
rect 198582 -14 198653 0
rect 198704 -14 198766 0
rect 198785 -14 198858 0
rect 198980 -14 199042 0
rect 199339 -14 199410 0
rect 199707 -14 199778 0
rect 200234 -14 200299 0
rect 200443 -14 200514 0
rect 201039 -14 201112 0
rect 201363 -14 201434 0
rect 201618 -14 201680 0
rect 201922 -14 202037 0
rect 202262 -14 202324 0
rect 202467 -14 202538 0
rect 202559 -14 202630 0
rect 202743 -14 202814 0
rect 202835 -14 202998 0
rect 203019 -14 203090 0
rect 203091 -14 203244 0
rect 203387 -14 203458 0
rect 203670 -14 203805 0
rect 203856 -14 203969 0
rect 204194 -14 204259 0
rect 204286 -14 204348 0
rect 204491 -14 204562 0
rect 204700 -14 204751 0
rect 204838 -14 204889 0
rect 205022 -14 205084 0
rect 205227 -14 205339 0
rect 205390 -14 205455 0
rect 205666 -14 205728 0
rect 206034 -14 206096 0
rect 206494 -14 206556 0
rect 206616 -14 206678 0
rect 206770 -14 206821 0
rect 207159 -14 207230 0
rect 207506 -14 207568 0
rect 207782 -14 207844 0
rect 208364 -14 208426 0
rect 208907 -14 208978 0
rect 209008 -14 209070 0
rect 209376 -14 209500 0
rect 209622 -14 209714 0
rect 209990 -14 210041 0
rect 210756 -14 210879 0
rect 211207 -14 211329 0
rect 211667 -14 211738 0
rect 212198 -14 212269 0
rect 212311 -14 212382 0
rect 212520 -14 212571 0
rect 212597 -14 212658 0
rect 212863 -14 212934 0
rect 212955 -14 213026 0
rect 213118 -14 213189 0
rect 213210 -14 213375 0
rect 215086 -14 215148 0
rect 215163 -14 215234 0
rect 215255 -14 215326 0
rect 215418 -14 215510 0
rect 215623 -14 215694 0
rect 215991 -14 216062 0
rect 216092 -14 216154 0
rect 216368 -14 216430 0
rect 216798 -14 216869 0
rect 216890 -14 216955 0
rect 217166 -14 217309 0
rect 217647 -14 217780 0
rect 217839 -14 217994 0
rect 218484 -14 218546 0
rect 218751 -14 218822 0
rect 220018 -14 220080 0
rect 220416 -14 220478 0
rect 220508 -14 220570 0
rect 220692 -14 220754 0
rect 220846 -14 220917 0
rect 220959 -14 221030 0
rect 221235 -14 221368 0
rect 221695 -14 221817 0
rect 222390 -14 222455 0
rect 222523 -14 222686 0
rect 222778 -14 223054 0
rect 224710 -14 224775 0
rect 224894 -14 225057 0
rect 225446 -14 225517 0
rect 226019 -14 226141 0
rect 226203 -14 226274 0
rect 226826 -14 226895 0
rect 227215 -14 227337 0
rect 227378 -14 227440 0
rect 228298 -14 228360 0
rect 228390 -14 228452 0
<< metal2 >>
rect 29642 0 29698 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 42522 0 42578 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 65706 0 65762 800
rect 66350 0 66406 800
rect 71502 0 71558 800
rect 72146 0 72202 800
rect 72790 0 72846 800
rect 73434 0 73490 800
<< obsm2 >>
rect 25124 25124 120832 218376
<< metal3 >>
rect 0 136008 800 136128
rect 0 135328 800 135448
rect 0 132608 800 132728
rect 230205 83648 231005 83768
rect 230205 80928 231005 81048
rect 230205 80248 231005 80368
rect 230205 78888 231005 79008
rect 230205 77528 231005 77648
<< obsm3 >>
rect 25000 0 226168 218376
rect 30782 -30 30886 0
rect 38566 -30 38686 0
rect 41470 -30 41538 0
rect 41630 -30 41708 0
rect 41814 -30 41890 0
rect 42758 -30 42854 0
rect 44098 -30 44214 0
rect 45218 -30 45290 0
rect 46966 -30 47046 0
rect 48958 -30 49082 0
rect 50140 -30 50218 0
rect 53282 -30 53406 0
rect 53573 -30 53651 0
rect 54340 -30 54418 0
rect 59584 -30 59662 0
rect 60013 -30 60091 0
rect 60410 -30 60534 0
rect 61502 -30 61580 0
rect 61778 -30 61856 0
rect 65918 -30 65996 0
rect 66304 -30 66382 0
rect 67266 -30 67390 0
rect 67482 -30 67594 0
rect 70486 -30 70610 0
rect 72280 -30 72358 0
rect 72830 -30 72910 0
rect 73830 -30 73908 0
rect 74270 -30 74382 0
rect 75224 -30 75380 0
rect 75776 -30 75854 0
rect 75900 -30 76004 0
rect 77202 -30 77326 0
rect 77340 -30 77418 0
rect 77478 -30 77602 0
rect 81558 -30 81636 0
rect 82093 -30 82171 0
rect 85758 -30 85882 0
rect 86704 -30 86782 0
rect 87245 -30 87323 0
rect 88426 -30 88550 0
rect 90588 -30 90666 0
rect 91140 -30 91218 0
rect 91462 -30 91586 0
rect 92198 -30 92414 0
rect 94070 -30 94148 0
rect 96830 -30 96908 0
rect 97488 -30 97644 0
rect 98408 -30 98532 0
rect 100478 -30 100602 0
rect 100878 -30 100998 0
rect 101730 -30 101968 0
rect 103376 -30 103500 0
rect 104558 -30 104678 0
rect 104986 -30 105110 0
rect 106938 -30 107042 0
rect 107686 -30 107870 0
rect 108114 -30 108316 0
rect 109020 -30 109098 0
rect 110138 -30 110262 0
rect 115014 -30 115138 0
rect 115690 -30 115768 0
rect 122130 -30 122208 0
rect 122328 -30 122452 0
rect 123556 -30 123634 0
rect 123740 -30 123818 0
rect 124062 -30 124140 0
rect 124260 -30 124338 0
rect 124352 -30 124430 0
rect 124582 -30 124706 0
rect 124812 -30 124890 0
rect 125718 -30 125822 0
rect 125870 -30 125948 0
rect 126054 -30 126132 0
rect 126192 -30 126348 0
rect 126454 -30 126532 0
rect 126652 -30 126730 0
rect 127770 -30 127834 0
rect 127986 -30 128110 0
rect 128584 -30 128662 0
rect 129122 -30 129306 0
rect 130828 -30 130916 0
rect 131252 -30 131330 0
rect 131574 -30 131698 0
rect 132080 -30 132158 0
rect 132894 -30 133002 0
rect 133092 -30 133262 0
rect 133860 -30 133980 0
rect 133998 -30 134182 0
rect 134918 -30 134996 0
rect 135254 -30 135332 0
rect 135484 -30 135562 0
rect 135576 -30 135654 0
rect 136022 -30 136100 0
rect 136128 -30 136284 0
rect 136312 -30 136468 0
rect 136496 -30 136574 0
rect 136588 -30 136744 0
rect 139578 -30 139702 0
rect 141266 -30 141380 0
rect 141924 -30 142080 0
rect 142338 -30 142462 0
rect 142936 -30 143092 0
rect 143452 -30 143566 0
rect 143796 -30 143874 0
rect 144270 -30 144394 0
rect 144960 -30 145038 0
rect 145222 -30 145300 0
rect 145420 -30 145682 0
rect 146110 -30 146234 0
rect 146340 -30 146418 0
rect 146478 -30 146694 0
rect 146850 -30 147048 0
rect 147218 -30 147338 0
rect 147858 -30 148074 0
rect 148414 -30 148534 0
rect 148732 -30 148810 0
rect 148916 -30 149086 0
rect 149270 -30 149348 0
rect 149426 -30 149546 0
rect 150020 -30 150098 0
rect 150296 -30 150374 0
rect 150604 -30 150682 0
rect 152214 -30 152292 0
rect 154160 -30 154238 0
rect 154560 -30 154698 0
rect 154804 -30 154960 0
rect 155172 -30 155250 0
rect 155954 -30 156078 0
rect 156492 -30 156630 0
rect 156690 -30 156906 0
rect 156920 -30 157090 0
rect 157748 -30 157904 0
rect 158378 -30 158456 0
rect 159666 -30 159744 0
rect 162794 -30 162872 0
rect 163176 -30 163254 0
rect 163692 -30 163806 0
rect 163820 -30 163898 0
rect 164050 -30 164266 0
rect 164330 -30 164450 0
rect 164832 -30 165034 0
rect 165462 -30 165540 0
rect 166212 -30 166290 0
rect 166906 -30 167026 0
rect 167946 -30 168024 0
rect 169188 -30 169266 0
rect 169418 -30 169602 0
rect 170352 -30 170508 0
rect 171364 -30 171442 0
rect 171456 -30 171612 0
rect 171732 -30 171810 0
rect 171916 -30 172072 0
rect 172698 -30 172822 0
rect 173622 -30 173926 0
rect 173940 -30 174018 0
rect 174110 -30 174202 0
rect 174216 -30 174386 0
rect 174400 -30 174570 0
rect 176516 -30 176672 0
rect 177068 -30 177224 0
rect 177252 -30 177408 0
rect 177804 -30 177882 0
rect 178020 -30 178098 0
rect 178218 -30 178342 0
rect 178356 -30 178512 0
rect 178908 -30 179064 0
rect 179124 -30 179202 0
rect 179920 -30 179998 0
rect 180090 -30 180228 0
rect 180242 -30 180366 0
rect 180380 -30 180664 0
rect 180748 -30 180826 0
rect 182358 -30 182560 0
rect 182680 -30 182836 0
rect 183834 -30 183954 0
rect 184244 -30 184322 0
rect 184520 -30 184598 0
rect 184846 -30 185090 0
rect 185302 -30 185426 0
rect 185532 -30 185610 0
rect 185716 -30 185964 0
rect 186176 -30 186378 0
rect 187514 -30 187634 0
rect 187786 -30 188080 0
rect 191926 -30 192142 0
rect 192846 -30 192970 0
rect 193122 -30 193246 0
rect 193398 -30 193614 0
rect 193766 -30 193890 0
rect 193996 -30 194152 0
rect 194824 -30 194902 0
rect 195008 -30 195316 0
rect 195468 -30 195546 0
rect 196052 -30 196130 0
rect 196604 -30 196682 0
rect 196756 -30 196834 0
rect 197110 -30 197188 0
rect 197446 -30 197708 0
rect 197722 -30 198030 0
rect 198918 -30 199042 0
rect 200054 -30 200132 0
rect 200160 -30 200238 0
rect 201080 -30 201158 0
rect 201908 -30 202078 0
rect 202322 -30 202538 0
rect 202598 -30 202722 0
rect 202966 -30 203274 0
rect 203430 -30 203664 0
rect 203918 -30 203996 0
rect 204208 -30 204286 0
rect 204442 -30 204562 0
rect 204700 -30 204838 0
rect 206048 -30 206126 0
rect 206646 -30 206848 0
rect 208072 -30 208150 0
rect 208854 -30 208978 0
rect 210422 -30 210542 0
rect 211370 -30 211448 0
rect 212396 -30 212658 0
rect 213210 -30 213394 0
rect 213762 -30 213840 0
rect 213914 -30 214038 0
rect 214558 -30 214682 0
rect 214880 -30 215036 0
rect 215602 -30 215680 0
rect 217028 -30 217106 0
rect 219070 -30 219268 0
rect 221274 -30 221398 0
rect 221738 -30 221858 0
rect 222778 -30 222962 0
rect 223528 -30 223698 0
rect 224494 -30 224618 0
rect 224816 -30 225064 0
rect 225354 -30 225432 0
rect 225506 -30 225630 0
rect 225966 -30 226168 0
<< metal4 >>
rect -3716 -2644 -3396 235476
rect -3056 -1984 -2736 234816
rect -2396 -1324 -2076 234156
rect -1736 -664 -1416 233496
rect -1076 -4 -756 232836
rect -416 656 -96 232176
rect 4208 -2644 4528 235476
rect 4868 -2644 5188 235476
rect 5528 -2644 5848 235476
rect 6188 -2644 6508 235476
rect 6848 -2644 7168 235476
rect 7508 -2644 7828 235476
rect 34928 218496 35248 235476
rect 35588 218496 35908 235476
rect 36248 218496 36568 235476
rect 36908 218496 37228 235476
rect 37568 218620 37888 235476
rect 38228 218620 38548 235476
rect 65648 218620 65968 235476
rect 66308 218620 66628 235476
rect 66968 218620 67288 235476
rect 67628 218620 67948 235476
rect 68288 218496 68608 235476
rect 68948 218620 69268 235476
rect 96368 218496 96688 235476
rect 97028 218620 97348 235476
rect 97688 218496 98008 235476
rect 98348 218620 98668 235476
rect 99008 218496 99328 235476
rect 99668 218620 99988 235476
rect 34928 104496 35248 139004
rect 35588 104496 35908 139004
rect 65648 104620 65968 139004
rect 66308 104496 66628 138880
rect 96368 104496 96688 139004
rect 97028 104496 97348 139004
rect 34928 -2644 35248 25004
rect 35588 -2644 35908 25004
rect 36248 -2644 36568 25004
rect 36908 -2644 37228 25004
rect 37568 -2644 37888 25004
rect 38228 -2644 38548 25004
rect 65648 -2644 65968 24880
rect 66308 -2644 66628 24880
rect 66968 -2644 67288 24880
rect 67628 -2644 67948 24880
rect 68288 -2644 68608 24880
rect 68948 -2644 69268 24880
rect 96368 -2644 96688 25004
rect 97028 -2644 97348 25004
rect 97688 -2644 98008 25004
rect 98348 -2644 98668 25004
rect 99008 -2644 99328 25004
rect 99668 -2644 99988 25004
rect 127088 -2644 127408 235476
rect 127748 -2644 128068 235476
rect 128408 -2644 128728 235476
rect 129068 -2644 129388 235476
rect 129728 -2644 130048 235476
rect 130388 -2644 130708 235476
rect 157808 -2644 158128 235476
rect 158468 -2644 158788 235476
rect 159128 -2644 159448 235476
rect 159788 -2644 160108 235476
rect 160448 -2644 160768 235476
rect 161108 -2644 161428 235476
rect 188528 -2644 188848 235476
rect 189188 -2644 189508 235476
rect 189848 -2644 190168 235476
rect 190508 -2644 190828 235476
rect 191168 -2644 191488 235476
rect 191828 -2644 192148 235476
rect 219248 -2644 219568 235476
rect 219908 -2644 220228 235476
rect 220568 -2644 220888 235476
rect 221228 -2644 221548 235476
rect 221888 -2644 222208 235476
rect 222548 -2644 222868 235476
rect 231016 656 231336 232176
rect 231676 -4 231996 232836
rect 232336 -664 232656 233496
rect 232996 -1324 233316 234156
rect 233656 -1984 233976 234816
rect 234316 -2644 234636 235476
<< obsm4 >>
rect 25124 218416 34848 218500
rect 35328 218416 35508 218500
rect 35988 218416 36168 218500
rect 36648 218416 36828 218500
rect 37308 218416 68208 218500
rect 68688 218416 96288 218500
rect 96768 218416 97608 218500
rect 98088 218416 98928 218500
rect 99408 218416 127008 218500
rect 25124 139084 127008 218416
rect 25124 104416 34848 139084
rect 35328 104416 35508 139084
rect 35988 104540 65568 139084
rect 66048 138960 96288 139084
rect 66048 104540 66228 138960
rect 35988 104416 66228 104540
rect 66708 104416 96288 138960
rect 96768 104416 96948 139084
rect 97428 104416 127008 139084
rect 25124 25084 127008 104416
rect 25124 0 34848 25084
rect 35328 0 35508 25084
rect 35988 0 36168 25084
rect 36648 0 36828 25084
rect 37308 0 37488 25084
rect 37968 0 38148 25084
rect 38628 24960 96288 25084
rect 38628 0 65568 24960
rect 66048 0 66228 24960
rect 66708 0 66888 24960
rect 67368 0 67548 24960
rect 68028 0 68208 24960
rect 68688 0 68868 24960
rect 69348 0 96288 24960
rect 96768 0 96948 25084
rect 97428 0 97608 25084
rect 98088 0 98268 25084
rect 98748 0 98928 25084
rect 99408 0 99588 25084
rect 100068 0 127008 25084
rect 126102 -124 126162 0
rect 126700 -124 126760 0
rect 127488 0 127668 218500
rect 128148 0 128328 218500
rect 128808 0 128988 218500
rect 129468 0 129648 218500
rect 130128 0 130308 218500
rect 130788 0 157728 218500
rect 135440 -124 135500 0
rect 145652 -124 145712 0
rect 149516 -124 149576 0
rect 154208 -124 154268 0
rect 157060 -124 157120 0
rect 158208 0 158388 218500
rect 158868 0 159048 218500
rect 159528 0 159708 218500
rect 160188 0 160368 218500
rect 160848 0 161028 218500
rect 161508 0 188448 218500
rect 164420 -124 164480 0
rect 171504 -124 171564 0
rect 171964 -124 172024 0
rect 172470 -124 172530 0
rect 172792 -124 172852 0
rect 176564 -124 176624 0
rect 177852 -124 177912 0
rect 177944 -124 178004 0
rect 178404 -124 178464 0
rect 180198 -124 180258 0
rect 180336 -124 180396 0
rect 182452 -124 182512 0
rect 182728 -124 182788 0
rect 183740 -124 183800 0
rect 188928 0 189108 218500
rect 189588 0 189768 218500
rect 190248 0 190428 218500
rect 190908 0 191088 218500
rect 191568 0 191748 218500
rect 192228 0 219168 218500
rect 202508 -124 202568 0
rect 203060 -124 203120 0
rect 206096 -124 206156 0
rect 219648 0 219828 218500
rect 220308 0 220488 218500
rect 220968 0 221148 218500
rect 221628 0 221808 218500
rect 222288 0 222468 218500
rect 222948 0 224924 218500
rect 224864 -124 224924 0
<< metal5 >>
rect -3716 235156 234636 235476
rect -3056 234496 233976 234816
rect -2396 233836 233316 234156
rect -1736 233176 232656 233496
rect -1076 232516 231996 232836
rect -416 231856 231336 232176
rect -3716 223098 234636 223418
rect -3716 222438 234636 222758
rect -3716 221778 234636 222098
rect -3716 221118 234636 221438
rect -3716 220458 234636 220778
rect -3716 219798 234636 220118
rect -3716 192462 234636 192782
rect -3716 191802 234636 192122
rect -3716 191142 234636 191462
rect -3716 190482 234636 190802
rect -3716 189822 234636 190142
rect -3716 189162 234636 189482
rect -3716 161826 234636 162146
rect -3716 161166 234636 161486
rect -3716 160506 234636 160826
rect -3716 159846 234636 160166
rect -3716 159186 234636 159506
rect -3716 158526 234636 158846
rect -3716 131190 234636 131510
rect -3716 130530 234636 130850
rect -3716 129870 234636 130190
rect -3716 129210 234636 129530
rect -3716 128550 234636 128870
rect -3716 127890 234636 128210
rect -3716 100554 234636 100874
rect -3716 99894 234636 100214
rect -3716 99234 234636 99554
rect -3716 98574 234636 98894
rect -3716 97914 234636 98234
rect -3716 97254 234636 97574
rect -3716 69918 234636 70238
rect -3716 69258 234636 69578
rect -3716 68598 234636 68918
rect -3716 67938 234636 68258
rect -3716 67278 234636 67598
rect -3716 66618 234636 66938
rect -3716 39282 234636 39602
rect -3716 38622 234636 38942
rect -3716 37962 234636 38282
rect -3716 37302 234636 37622
rect -3716 36642 234636 36962
rect -3716 35982 234636 36302
rect -3716 8646 234636 8966
rect -3716 7986 234636 8306
rect -3716 7326 234636 7646
rect -3716 6666 234636 6986
rect -3716 6006 234636 6326
rect -3716 5346 234636 5666
rect -416 656 231336 976
rect -1076 -4 231996 316
rect -1736 -664 232656 -344
rect -2396 -1324 233316 -1004
rect -3056 -1984 233976 -1664
rect -3716 -2644 234636 -2324
<< labels >>
rlabel metal4 s -2396 -1324 -2076 234156 4 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2396 -1324 233316 -1004 8 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2396 233836 233316 234156 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 232996 -1324 233316 234156 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6188 -2644 6508 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 36908 -2644 37228 25004 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 36908 218496 37228 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67628 -2644 67948 24880 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 67628 218620 67948 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98348 -2644 98668 25004 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98348 218620 98668 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 129068 -2644 129388 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 159788 -2644 160108 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 190508 -2644 190828 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 221228 -2644 221548 235476 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 7326 234636 7646 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 37962 234636 38282 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 68598 234636 68918 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 99234 234636 99554 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 129870 234636 130190 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 160506 234636 160826 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 191142 234636 191462 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -3716 221778 234636 222098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s -3716 -2644 -3396 235476 4 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 -2644 234636 -2324 8 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 235156 234636 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 234316 -2644 234636 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 7508 -2644 7828 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 38228 -2644 38548 25004 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 38228 218620 38548 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 68948 -2644 69268 24880 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 68948 218620 69268 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 99668 -2644 99988 25004 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 99668 218620 99988 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 130388 -2644 130708 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 161108 -2644 161428 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 191828 -2644 192148 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s 222548 -2644 222868 235476 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 8646 234636 8966 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 39282 234636 39602 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 69918 234636 70238 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 100554 234636 100874 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 131190 234636 131510 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 161826 234636 162146 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 192462 234636 192782 6 VNB
port 2 nsew ground bidirectional
rlabel metal5 s -3716 223098 234636 223418 6 VNB
port 2 nsew ground bidirectional
rlabel metal4 s -3056 -1984 -2736 234816 4 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3056 -1984 233976 -1664 8 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3056 234496 233976 234816 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 233656 -1984 233976 234816 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 6848 -2644 7168 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 37568 -2644 37888 25004 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 37568 218620 37888 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 68288 -2644 68608 24880 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 68288 218496 68608 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 99008 -2644 99328 25004 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 99008 218496 99328 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 129728 -2644 130048 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 160448 -2644 160768 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 191168 -2644 191488 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s 221888 -2644 222208 235476 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 7986 234636 8306 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 38622 234636 38942 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 69258 234636 69578 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 99894 234636 100214 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 130530 234636 130850 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 161166 234636 161486 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 191802 234636 192122 6 VPB
port 3 nsew power bidirectional
rlabel metal5 s -3716 222438 234636 222758 6 VPB
port 3 nsew power bidirectional
rlabel metal4 s -1736 -664 -1416 233496 4 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -1736 -664 232656 -344 8 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -1736 233176 232656 233496 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 232336 -664 232656 233496 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 5528 -2644 5848 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 36248 -2644 36568 25004 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 36248 218496 36568 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 66968 -2644 67288 24880 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 66968 218620 67288 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 97688 -2644 98008 25004 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 97688 218496 98008 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 128408 -2644 128728 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 159128 -2644 159448 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 189848 -2644 190168 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 220568 -2644 220888 235476 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 6666 234636 6986 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 37302 234636 37622 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 67938 234636 68258 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 98574 234636 98894 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 129210 234636 129530 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 159846 234636 160166 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 190482 234636 190802 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s -3716 221118 234636 221438 6 VPWR
port 4 nsew power bidirectional
rlabel metal2 s 29642 0 29698 800 6 clk
port 5 nsew signal input
rlabel metal3 s 230205 77528 231005 77648 6 input_gpio_pins[0]
port 6 nsew signal input
rlabel metal3 s 230205 78888 231005 79008 6 input_gpio_pins[1]
port 7 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 instructions[0]
port 8 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 instructions[1]
port 9 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 instructions[2]
port 10 nsew signal output
rlabel metal3 s 230205 80928 231005 81048 6 output_gpio_pins[0]
port 11 nsew signal output
rlabel metal3 s 230205 80248 231005 80368 6 output_gpio_pins[1]
port 12 nsew signal output
rlabel metal3 s 230205 83648 231005 83768 6 output_gpio_pins[2]
port 13 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 resetn
port 14 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 uart_rx_break
port 15 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 uart_rx_data[0]
port 16 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 uart_rx_data[1]
port 17 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 uart_rx_data[2]
port 18 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 uart_rx_data[3]
port 19 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 uart_rx_data[4]
port 20 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 uart_rx_data[5]
port 21 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 uart_rx_data[6]
port 22 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 uart_rx_data[7]
port 23 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 uart_rx_en
port 24 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 uart_rx_valid
port 25 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 uart_rxd
port 26 nsew signal input
rlabel metal4 s -416 656 -96 232176 4 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -416 656 231336 976 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -416 231856 231336 232176 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 231016 656 231336 232176 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 4208 -2644 4528 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 34928 -2644 35248 25004 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 34928 104496 35248 139004 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 34928 218496 35248 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 65648 -2644 65968 24880 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 65648 104620 65968 139004 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 65648 218620 65968 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 96368 -2644 96688 25004 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 96368 104496 96688 139004 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 96368 218496 96688 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 127088 -2644 127408 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 157808 -2644 158128 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 188528 -2644 188848 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 219248 -2644 219568 235476 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 5346 234636 5666 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 35982 234636 36302 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 66618 234636 66938 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 97254 234636 97574 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 127890 234636 128210 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 158526 234636 158846 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 189162 234636 189482 6 vccd1
port 27 nsew power bidirectional
rlabel metal5 s -3716 219798 234636 220118 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s -1076 -4 -756 232836 4 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -1076 -4 231996 316 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -1076 232516 231996 232836 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 231676 -4 231996 232836 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 4868 -2644 5188 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 35588 -2644 35908 25004 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 35588 104496 35908 139004 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 35588 218496 35908 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 66308 -2644 66628 24880 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 66308 104496 66628 138880 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 66308 218620 66628 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 97028 -2644 97348 25004 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 97028 104496 97348 139004 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 97028 218620 97348 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 127748 -2644 128068 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 158468 -2644 158788 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 189188 -2644 189508 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 219908 -2644 220228 235476 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 6006 234636 6326 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 36642 234636 36962 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 67278 234636 67598 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 97914 234636 98234 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 128550 234636 128870 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 159186 234636 159506 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 189822 234636 190142 6 vssd1
port 28 nsew ground bidirectional
rlabel metal5 s -3716 220458 234636 220778 6 vssd1
port 28 nsew ground bidirectional
rlabel metal2 s 46386 0 46442 800 6 write_done
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 231005 233149
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21935044
string GDS_FILE /openlane/designs/kanish/runs/RUN_2023.11.14_19.09.44/results/signoff/wrapper.magic.gds
string GDS_START 10660972
<< end >>

